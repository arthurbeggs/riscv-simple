module scan2ascii (
	input wire [7:0] scan,
	input wire shift,
	output wire [7:0] ascii
);

wire [1024:0] sem_shift;
wire [1024:0] com_shift;

wire  [10:0] indice = scan < 8'h80 ? 11'd1023 - (scan << 3) : 11'b0;

assign ascii = shift ? com_shift[ indice -: 8 ] : sem_shift[ indice -: 8 ];


assign sem_shift = {
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h71, 8'h31, 8'h00, 8'h00, 8'h00, 8'h7a, 8'h73, 8'h61, 8'h77, 8'h32, 8'h00,  
	8'h00, 8'h63, 8'h78, 8'h64, 8'h65, 8'h34, 8'h33, 8'h00, 8'h00, 8'h20, 8'h76, 8'h66, 8'h74, 8'h72, 8'h35, 8'h00, 
	8'h00, 8'h6e, 8'h62, 8'h68, 8'h67, 8'h79, 8'h36, 8'h00, 8'h00, 8'h00, 8'h6d, 8'h6a, 8'h75, 8'h37, 8'h38, 8'h00, 
	8'h00, 8'h2c, 8'h6b, 8'h69, 8'h6f, 8'h30, 8'h39, 8'h00, 8'h00, 8'h2e, 8'h2f, 8'h6c, 8'h3b, 8'h70, 8'h2d, 8'h00,  
	8'h00, 8'h00, 8'h27, 8'h00, 8'h00, 8'h3d, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h5b, 8'h00, 8'h5d, 8'h00, 8'h00, 
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h00, 8'h34, 8'h37, 8'h00, 8'h00, 8'h00,  
	8'h30, 8'h2e, 8'h32, 8'h35, 8'h36, 8'h38, 8'h00, 8'h00, 8'h00, 8'h2b, 8'h33, 8'h2d, 8'h2a, 8'h39, 8'h00, 8'h00
	};
	
assign com_shift = {
   8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h21, 8'h00, 8'h00, 8'h00, 8'h5a, 8'h53, 8'h41, 8'h57, 8'h40, 8'h00, 
	8'h00, 8'h43, 8'h58, 8'h44, 8'h45, 8'h24, 8'h23, 8'h00, 8'h00, 8'h00, 8'h56, 8'h46, 8'h54, 8'h52, 8'h25, 8'h00, 
	8'h00, 8'h4e, 8'h42, 8'h48, 8'h47, 8'h59, 8'h5e, 8'h00, 8'h00, 8'h00, 8'h4d, 8'h4a, 8'h55, 8'h26, 8'h2a, 8'h00, 
	8'h00, 8'h3c, 8'h4b, 8'h49, 8'h4f, 8'h29, 8'h28, 8'h00, 8'h00, 8'h3e, 8'h3f, 8'h4c, 8'h3a, 8'h50, 8'h5f, 8'h00, 
	8'h00, 8'h00, 8'h22, 8'h00, 8'h00, 8'h2b, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7b, 8'h00, 8'h7d, 8'h00, 8'h00, 
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 
	8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00	
	};


endmodule
	